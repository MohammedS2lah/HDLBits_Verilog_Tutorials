* Step one
---------------
module top_module( output one );

// Insert your code here
    assign one = 1'b1;

endmodule


----------------

* Zero
----------------
module top_module(
    output zero
);// Module body starts after semicolon
	assign zero = 1'b0;
endmodule
